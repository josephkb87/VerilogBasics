// Combinational logic vs Sequential logic